`timescale 1ns/1ns





module processor(input clk);

wire clk;



endmodule

